`timescale 1ns/1ps
module sample ();
  $display("This is a sample code");
endmodule
